
module dikkekoek (
	clk_clk,
	reset_reset_n,
	camera_input_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	input	[11:0]	camera_input_external_connection_export;
endmodule
