
module camerametnios (
	camera_input_0_external_connection_export,
	camera_input_1_external_connection_export,
	camera_input_2_external_connection_export,
	camera_input_3_external_connection_export,
	camera_input_4_external_connection_export,
	camera_input_5_external_connection_export,
	camera_input_6_external_connection_export,
	camera_input_7_external_connection_export,
	camera_input_8_external_connection_export,
	camera_input_9_external_connection_export,
	clk_clk,
	reset_reset_n);	

	input	[14:0]	camera_input_0_external_connection_export;
	input	[14:0]	camera_input_1_external_connection_export;
	input	[14:0]	camera_input_2_external_connection_export;
	input	[14:0]	camera_input_3_external_connection_export;
	input	[14:0]	camera_input_4_external_connection_export;
	input	[14:0]	camera_input_5_external_connection_export;
	input	[14:0]	camera_input_6_external_connection_export;
	input	[14:0]	camera_input_7_external_connection_export;
	input	[14:0]	camera_input_8_external_connection_export;
	input	[14:0]	camera_input_9_external_connection_export;
	input		clk_clk;
	input		reset_reset_n;
endmodule
