-- nios_system.vhd

-- Generated using ACDS version 16.1 203

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_system is
	port (
		cam_in_0_external_connection_export : in    std_logic_vector(14 downto 0) := (others => '0'); -- cam_in_0_external_connection.export
		cam_in_1_external_connection_export : in    std_logic_vector(14 downto 0) := (others => '0'); -- cam_in_1_external_connection.export
		cam_in_2_external_connection_export : in    std_logic_vector(14 downto 0) := (others => '0'); -- cam_in_2_external_connection.export
		cam_in_3_external_connection_export : in    std_logic_vector(14 downto 0) := (others => '0'); -- cam_in_3_external_connection.export
		cam_in_4_external_connection_export : in    std_logic_vector(14 downto 0) := (others => '0'); -- cam_in_4_external_connection.export
		cam_in_5_external_connection_export : in    std_logic_vector(14 downto 0) := (others => '0'); -- cam_in_5_external_connection.export
		cam_in_6_external_connection_export : in    std_logic_vector(14 downto 0) := (others => '0'); -- cam_in_6_external_connection.export
		cam_in_7_external_connection_export : in    std_logic_vector(14 downto 0) := (others => '0'); -- cam_in_7_external_connection.export
		cam_in_8_external_connection_export : in    std_logic_vector(14 downto 0) := (others => '0'); -- cam_in_8_external_connection.export
		cam_in_9_external_connection_export : in    std_logic_vector(14 downto 0) := (others => '0'); -- cam_in_9_external_connection.export
		flash_ADDR                          : out   std_logic_vector(22 downto 0);                    --                        flash.ADDR
		flash_CE_N                          : out   std_logic;                                        --                             .CE_N
		flash_OE_N                          : out   std_logic;                                        --                             .OE_N
		flash_WE_N                          : out   std_logic;                                        --                             .WE_N
		flash_RST_N                         : out   std_logic;                                        --                             .RST_N
		flash_DQ                            : inout std_logic_vector(7 downto 0)  := (others => '0'); --                             .DQ
		sdram_addr                          : out   std_logic_vector(12 downto 0);                    --                        sdram.addr
		sdram_ba                            : out   std_logic_vector(1 downto 0);                     --                             .ba
		sdram_cas_n                         : out   std_logic;                                        --                             .cas_n
		sdram_cke                           : out   std_logic;                                        --                             .cke
		sdram_cs_n                          : out   std_logic;                                        --                             .cs_n
		sdram_dq                            : inout std_logic_vector(31 downto 0) := (others => '0'); --                             .dq
		sdram_dqm                           : out   std_logic_vector(3 downto 0);                     --                             .dqm
		sdram_ras_n                         : out   std_logic;                                        --                             .ras_n
		sdram_we_n                          : out   std_logic;                                        --                             .we_n
		sdram_clk_clk                       : out   std_logic;                                        --                    sdram_clk.clk
		sram_DQ                             : inout std_logic_vector(15 downto 0) := (others => '0'); --                         sram.DQ
		sram_ADDR                           : out   std_logic_vector(19 downto 0);                    --                             .ADDR
		sram_LB_N                           : out   std_logic;                                        --                             .LB_N
		sram_UB_N                           : out   std_logic;                                        --                             .UB_N
		sram_CE_N                           : out   std_logic;                                        --                             .CE_N
		sram_OE_N                           : out   std_logic;                                        --                             .OE_N
		sram_WE_N                           : out   std_logic;                                        --                             .WE_N
		system_pll_ref_clk_clk              : in    std_logic                     := '0';             --           system_pll_ref_clk.clk
		system_pll_ref_reset_reset          : in    std_logic                     := '0'              --         system_pll_ref_reset.reset
	);
end entity nios_system;

architecture rtl of nios_system is
	component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface is
		generic (
			FLASH_MEMORY_ADDRESS_WIDTH : integer := 22
		);
		port (
			i_avalon_chip_select       : in    std_logic                     := 'X';             -- chipselect
			i_avalon_write             : in    std_logic                     := 'X';             -- write
			i_avalon_read              : in    std_logic                     := 'X';             -- read
			i_avalon_address           : in    std_logic_vector(20 downto 0) := (others => 'X'); -- address
			i_avalon_byteenable        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			i_avalon_writedata         : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			o_avalon_readdata          : out   std_logic_vector(31 downto 0);                    -- readdata
			o_avalon_waitrequest       : out   std_logic;                                        -- waitrequest
			i_clock                    : in    std_logic                     := 'X';             -- clk
			i_reset_n                  : in    std_logic                     := 'X';             -- reset_n
			FL_ADDR                    : out   std_logic_vector(22 downto 0);                    -- export
			FL_CE_N                    : out   std_logic;                                        -- export
			FL_OE_N                    : out   std_logic;                                        -- export
			FL_WE_N                    : out   std_logic;                                        -- export
			FL_RST_N                   : out   std_logic;                                        -- export
			FL_DQ                      : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			i_avalon_erase_write       : in    std_logic                     := 'X';             -- write
			i_avalon_erase_read        : in    std_logic                     := 'X';             -- read
			i_avalon_erase_byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			i_avalon_erase_writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			i_avalon_erase_chip_select : in    std_logic                     := 'X';             -- chipselect
			o_avalon_erase_readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			o_avalon_erase_waitrequest : out   std_logic                                         -- waitrequest
		);
	end component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface;

	component nios_system_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_system_JTAG_UART;

	component nios_system_Nios2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			d_address                           : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios_system_Nios2;

	component nios_system_Nios2_2nd_Core is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			d_address                           : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios_system_Nios2_2nd_Core;

	component nios_system_SDRAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component nios_system_SDRAM;

	component nios_system_SRAM is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component nios_system_SRAM;

	component nios_system_System_PLL is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component nios_system_System_PLL;

	component nios_system_cam_in_0 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(14 downto 0) := (others => 'X')  -- export
		);
	end component nios_system_cam_in_0;

	component nios_system_mm_interconnect_0 is
		port (
			System_PLL_sys_clk_clk                           : in  std_logic                     := 'X';             -- clk
			cam_in_8_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			JTAG_UART_reset_reset_bridge_in_reset_reset      : in  std_logic                     := 'X';             -- reset
			Nios2_2nd_Core_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Nios2_reset_reset_bridge_in_reset_reset          : in  std_logic                     := 'X';             -- reset
			Nios2_data_master_address                        : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			Nios2_data_master_waitrequest                    : out std_logic;                                        -- waitrequest
			Nios2_data_master_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Nios2_data_master_read                           : in  std_logic                     := 'X';             -- read
			Nios2_data_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			Nios2_data_master_write                          : in  std_logic                     := 'X';             -- write
			Nios2_data_master_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Nios2_data_master_debugaccess                    : in  std_logic                     := 'X';             -- debugaccess
			Nios2_instruction_master_address                 : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			Nios2_instruction_master_waitrequest             : out std_logic;                                        -- waitrequest
			Nios2_instruction_master_read                    : in  std_logic                     := 'X';             -- read
			Nios2_instruction_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			Nios2_instruction_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			Nios2_2nd_Core_data_master_address               : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			Nios2_2nd_Core_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			Nios2_2nd_Core_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Nios2_2nd_Core_data_master_read                  : in  std_logic                     := 'X';             -- read
			Nios2_2nd_Core_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			Nios2_2nd_Core_data_master_write                 : in  std_logic                     := 'X';             -- write
			Nios2_2nd_Core_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Nios2_2nd_Core_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			Nios2_2nd_Core_instruction_master_address        : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			Nios2_2nd_Core_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			Nios2_2nd_Core_instruction_master_read           : in  std_logic                     := 'X';             -- read
			Nios2_2nd_Core_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			Nios2_2nd_Core_instruction_master_readdatavalid  : out std_logic;                                        -- readdatavalid
			cam_in_0_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			cam_in_0_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cam_in_1_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			cam_in_1_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cam_in_2_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			cam_in_2_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cam_in_3_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			cam_in_3_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cam_in_4_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			cam_in_4_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cam_in_5_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			cam_in_5_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cam_in_6_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			cam_in_6_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cam_in_7_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			cam_in_7_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cam_in_8_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			cam_in_8_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cam_in_9_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			cam_in_9_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Flash_flash_data_address                         : out std_logic_vector(20 downto 0);                    -- address
			Flash_flash_data_write                           : out std_logic;                                        -- write
			Flash_flash_data_read                            : out std_logic;                                        -- read
			Flash_flash_data_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Flash_flash_data_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			Flash_flash_data_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			Flash_flash_data_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			Flash_flash_data_chipselect                      : out std_logic;                                        -- chipselect
			Flash_flash_erase_control_write                  : out std_logic;                                        -- write
			Flash_flash_erase_control_read                   : out std_logic;                                        -- read
			Flash_flash_erase_control_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Flash_flash_erase_control_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			Flash_flash_erase_control_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			Flash_flash_erase_control_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			Flash_flash_erase_control_chipselect             : out std_logic;                                        -- chipselect
			JTAG_UART_avalon_jtag_slave_address              : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_avalon_jtag_slave_write                : out std_logic;                                        -- write
			JTAG_UART_avalon_jtag_slave_read                 : out std_logic;                                        -- read
			JTAG_UART_avalon_jtag_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_avalon_jtag_slave_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_avalon_jtag_slave_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect           : out std_logic;                                        -- chipselect
			JTAG_UART_2nd_Core_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_2nd_Core_avalon_jtag_slave_write       : out std_logic;                                        -- write
			JTAG_UART_2nd_Core_avalon_jtag_slave_read        : out std_logic;                                        -- read
			JTAG_UART_2nd_Core_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_2nd_Core_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_2nd_Core_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_2nd_Core_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			Nios2_debug_mem_slave_address                    : out std_logic_vector(8 downto 0);                     -- address
			Nios2_debug_mem_slave_write                      : out std_logic;                                        -- write
			Nios2_debug_mem_slave_read                       : out std_logic;                                        -- read
			Nios2_debug_mem_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Nios2_debug_mem_slave_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			Nios2_debug_mem_slave_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			Nios2_debug_mem_slave_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			Nios2_debug_mem_slave_debugaccess                : out std_logic;                                        -- debugaccess
			Nios2_2nd_Core_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			Nios2_2nd_Core_debug_mem_slave_write             : out std_logic;                                        -- write
			Nios2_2nd_Core_debug_mem_slave_read              : out std_logic;                                        -- read
			Nios2_2nd_Core_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Nios2_2nd_Core_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			Nios2_2nd_Core_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			Nios2_2nd_Core_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			Nios2_2nd_Core_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			SDRAM_s1_address                                 : out std_logic_vector(24 downto 0);                    -- address
			SDRAM_s1_write                                   : out std_logic;                                        -- write
			SDRAM_s1_read                                    : out std_logic;                                        -- read
			SDRAM_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SDRAM_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			SDRAM_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			SDRAM_s1_readdatavalid                           : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_s1_waitrequest                             : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_s1_chipselect                              : out std_logic;                                        -- chipselect
			SRAM_avalon_sram_slave_address                   : out std_logic_vector(19 downto 0);                    -- address
			SRAM_avalon_sram_slave_write                     : out std_logic;                                        -- write
			SRAM_avalon_sram_slave_read                      : out std_logic;                                        -- read
			SRAM_avalon_sram_slave_readdata                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SRAM_avalon_sram_slave_writedata                 : out std_logic_vector(15 downto 0);                    -- writedata
			SRAM_avalon_sram_slave_byteenable                : out std_logic_vector(1 downto 0);                     -- byteenable
			SRAM_avalon_sram_slave_readdatavalid             : in  std_logic                     := 'X'              -- readdatavalid
		);
	end component nios_system_mm_interconnect_0;

	component nios_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_system_irq_mapper;

	component nios_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_system_rst_controller;

	component nios_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_system_rst_controller_001;

	component nios_system_rst_controller_003 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_in2      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_system_rst_controller_003;

	signal system_pll_sys_clk_clk                                                 : std_logic;                     -- System_PLL:sys_clk_clk -> [Flash:i_clock, JTAG_UART:clk, JTAG_UART_2nd_Core:clk, Nios2:clk, Nios2_2nd_Core:clk, SDRAM:clk, SRAM:clk, cam_in_0:clk, cam_in_1:clk, cam_in_2:clk, cam_in_3:clk, cam_in_4:clk, cam_in_5:clk, cam_in_6:clk, cam_in_7:clk, cam_in_8:clk, cam_in_9:clk, irq_mapper:clk, irq_mapper_001:clk, mm_interconnect_0:System_PLL_sys_clk_clk, rst_controller:clk, rst_controller_001:clk, rst_controller_002:clk, rst_controller_003:clk]
	signal nios2_data_master_readdata                                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:Nios2_data_master_readdata -> Nios2:d_readdata
	signal nios2_data_master_waitrequest                                          : std_logic;                     -- mm_interconnect_0:Nios2_data_master_waitrequest -> Nios2:d_waitrequest
	signal nios2_data_master_debugaccess                                          : std_logic;                     -- Nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Nios2_data_master_debugaccess
	signal nios2_data_master_address                                              : std_logic_vector(28 downto 0); -- Nios2:d_address -> mm_interconnect_0:Nios2_data_master_address
	signal nios2_data_master_byteenable                                           : std_logic_vector(3 downto 0);  -- Nios2:d_byteenable -> mm_interconnect_0:Nios2_data_master_byteenable
	signal nios2_data_master_read                                                 : std_logic;                     -- Nios2:d_read -> mm_interconnect_0:Nios2_data_master_read
	signal nios2_data_master_write                                                : std_logic;                     -- Nios2:d_write -> mm_interconnect_0:Nios2_data_master_write
	signal nios2_data_master_writedata                                            : std_logic_vector(31 downto 0); -- Nios2:d_writedata -> mm_interconnect_0:Nios2_data_master_writedata
	signal nios2_2nd_core_data_master_readdata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:Nios2_2nd_Core_data_master_readdata -> Nios2_2nd_Core:d_readdata
	signal nios2_2nd_core_data_master_waitrequest                                 : std_logic;                     -- mm_interconnect_0:Nios2_2nd_Core_data_master_waitrequest -> Nios2_2nd_Core:d_waitrequest
	signal nios2_2nd_core_data_master_debugaccess                                 : std_logic;                     -- Nios2_2nd_Core:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Nios2_2nd_Core_data_master_debugaccess
	signal nios2_2nd_core_data_master_address                                     : std_logic_vector(28 downto 0); -- Nios2_2nd_Core:d_address -> mm_interconnect_0:Nios2_2nd_Core_data_master_address
	signal nios2_2nd_core_data_master_byteenable                                  : std_logic_vector(3 downto 0);  -- Nios2_2nd_Core:d_byteenable -> mm_interconnect_0:Nios2_2nd_Core_data_master_byteenable
	signal nios2_2nd_core_data_master_read                                        : std_logic;                     -- Nios2_2nd_Core:d_read -> mm_interconnect_0:Nios2_2nd_Core_data_master_read
	signal nios2_2nd_core_data_master_write                                       : std_logic;                     -- Nios2_2nd_Core:d_write -> mm_interconnect_0:Nios2_2nd_Core_data_master_write
	signal nios2_2nd_core_data_master_writedata                                   : std_logic_vector(31 downto 0); -- Nios2_2nd_Core:d_writedata -> mm_interconnect_0:Nios2_2nd_Core_data_master_writedata
	signal nios2_instruction_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Nios2_instruction_master_readdata -> Nios2:i_readdata
	signal nios2_instruction_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:Nios2_instruction_master_waitrequest -> Nios2:i_waitrequest
	signal nios2_instruction_master_address                                       : std_logic_vector(27 downto 0); -- Nios2:i_address -> mm_interconnect_0:Nios2_instruction_master_address
	signal nios2_instruction_master_read                                          : std_logic;                     -- Nios2:i_read -> mm_interconnect_0:Nios2_instruction_master_read
	signal nios2_instruction_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:Nios2_instruction_master_readdatavalid -> Nios2:i_readdatavalid
	signal nios2_2nd_core_instruction_master_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:Nios2_2nd_Core_instruction_master_readdata -> Nios2_2nd_Core:i_readdata
	signal nios2_2nd_core_instruction_master_waitrequest                          : std_logic;                     -- mm_interconnect_0:Nios2_2nd_Core_instruction_master_waitrequest -> Nios2_2nd_Core:i_waitrequest
	signal nios2_2nd_core_instruction_master_address                              : std_logic_vector(27 downto 0); -- Nios2_2nd_Core:i_address -> mm_interconnect_0:Nios2_2nd_Core_instruction_master_address
	signal nios2_2nd_core_instruction_master_read                                 : std_logic;                     -- Nios2_2nd_Core:i_read -> mm_interconnect_0:Nios2_2nd_Core_instruction_master_read
	signal nios2_2nd_core_instruction_master_readdatavalid                        : std_logic;                     -- mm_interconnect_0:Nios2_2nd_Core_instruction_master_readdatavalid -> Nios2_2nd_Core:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect               : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                 : std_logic_vector(31 downto 0); -- JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest              : std_logic;                     -- JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                     : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                    : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	signal mm_interconnect_0_sram_avalon_sram_slave_readdata                      : std_logic_vector(15 downto 0); -- SRAM:readdata -> mm_interconnect_0:SRAM_avalon_sram_slave_readdata
	signal mm_interconnect_0_sram_avalon_sram_slave_address                       : std_logic_vector(19 downto 0); -- mm_interconnect_0:SRAM_avalon_sram_slave_address -> SRAM:address
	signal mm_interconnect_0_sram_avalon_sram_slave_read                          : std_logic;                     -- mm_interconnect_0:SRAM_avalon_sram_slave_read -> SRAM:read
	signal mm_interconnect_0_sram_avalon_sram_slave_byteenable                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SRAM_avalon_sram_slave_byteenable -> SRAM:byteenable
	signal mm_interconnect_0_sram_avalon_sram_slave_readdatavalid                 : std_logic;                     -- SRAM:readdatavalid -> mm_interconnect_0:SRAM_avalon_sram_slave_readdatavalid
	signal mm_interconnect_0_sram_avalon_sram_slave_write                         : std_logic;                     -- mm_interconnect_0:SRAM_avalon_sram_slave_write -> SRAM:write
	signal mm_interconnect_0_sram_avalon_sram_slave_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:SRAM_avalon_sram_slave_writedata -> SRAM:writedata
	signal mm_interconnect_0_nios2_debug_mem_slave_readdata                       : std_logic_vector(31 downto 0); -- Nios2:debug_mem_slave_readdata -> mm_interconnect_0:Nios2_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_debug_mem_slave_waitrequest                    : std_logic;                     -- Nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:Nios2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_debug_mem_slave_debugaccess                    : std_logic;                     -- mm_interconnect_0:Nios2_debug_mem_slave_debugaccess -> Nios2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_debug_mem_slave_address                        : std_logic_vector(8 downto 0);  -- mm_interconnect_0:Nios2_debug_mem_slave_address -> Nios2:debug_mem_slave_address
	signal mm_interconnect_0_nios2_debug_mem_slave_read                           : std_logic;                     -- mm_interconnect_0:Nios2_debug_mem_slave_read -> Nios2:debug_mem_slave_read
	signal mm_interconnect_0_nios2_debug_mem_slave_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Nios2_debug_mem_slave_byteenable -> Nios2:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_debug_mem_slave_write                          : std_logic;                     -- mm_interconnect_0:Nios2_debug_mem_slave_write -> Nios2:debug_mem_slave_write
	signal mm_interconnect_0_nios2_debug_mem_slave_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Nios2_debug_mem_slave_writedata -> Nios2:debug_mem_slave_writedata
	signal mm_interconnect_0_flash_flash_data_chipselect                          : std_logic;                     -- mm_interconnect_0:Flash_flash_data_chipselect -> Flash:i_avalon_chip_select
	signal mm_interconnect_0_flash_flash_data_readdata                            : std_logic_vector(31 downto 0); -- Flash:o_avalon_readdata -> mm_interconnect_0:Flash_flash_data_readdata
	signal mm_interconnect_0_flash_flash_data_waitrequest                         : std_logic;                     -- Flash:o_avalon_waitrequest -> mm_interconnect_0:Flash_flash_data_waitrequest
	signal mm_interconnect_0_flash_flash_data_address                             : std_logic_vector(20 downto 0); -- mm_interconnect_0:Flash_flash_data_address -> Flash:i_avalon_address
	signal mm_interconnect_0_flash_flash_data_read                                : std_logic;                     -- mm_interconnect_0:Flash_flash_data_read -> Flash:i_avalon_read
	signal mm_interconnect_0_flash_flash_data_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Flash_flash_data_byteenable -> Flash:i_avalon_byteenable
	signal mm_interconnect_0_flash_flash_data_write                               : std_logic;                     -- mm_interconnect_0:Flash_flash_data_write -> Flash:i_avalon_write
	signal mm_interconnect_0_flash_flash_data_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:Flash_flash_data_writedata -> Flash:i_avalon_writedata
	signal mm_interconnect_0_flash_flash_erase_control_chipselect                 : std_logic;                     -- mm_interconnect_0:Flash_flash_erase_control_chipselect -> Flash:i_avalon_erase_chip_select
	signal mm_interconnect_0_flash_flash_erase_control_readdata                   : std_logic_vector(31 downto 0); -- Flash:o_avalon_erase_readdata -> mm_interconnect_0:Flash_flash_erase_control_readdata
	signal mm_interconnect_0_flash_flash_erase_control_waitrequest                : std_logic;                     -- Flash:o_avalon_erase_waitrequest -> mm_interconnect_0:Flash_flash_erase_control_waitrequest
	signal mm_interconnect_0_flash_flash_erase_control_read                       : std_logic;                     -- mm_interconnect_0:Flash_flash_erase_control_read -> Flash:i_avalon_erase_read
	signal mm_interconnect_0_flash_flash_erase_control_byteenable                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Flash_flash_erase_control_byteenable -> Flash:i_avalon_erase_byteenable
	signal mm_interconnect_0_flash_flash_erase_control_write                      : std_logic;                     -- mm_interconnect_0:Flash_flash_erase_control_write -> Flash:i_avalon_erase_write
	signal mm_interconnect_0_flash_flash_erase_control_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:Flash_flash_erase_control_writedata -> Flash:i_avalon_erase_writedata
	signal mm_interconnect_0_sdram_s1_chipselect                                  : std_logic;                     -- mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                    : std_logic_vector(31 downto 0); -- SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                 : std_logic;                     -- SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                     : std_logic_vector(24 downto 0); -- mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	signal mm_interconnect_0_sdram_s1_read                                        : std_logic;                     -- mm_interconnect_0:SDRAM_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SDRAM_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                               : std_logic;                     -- SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                       : std_logic;                     -- mm_interconnect_0:SDRAM_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	signal mm_interconnect_0_cam_in_8_s1_readdata                                 : std_logic_vector(31 downto 0); -- cam_in_8:readdata -> mm_interconnect_0:cam_in_8_s1_readdata
	signal mm_interconnect_0_cam_in_8_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:cam_in_8_s1_address -> cam_in_8:address
	signal mm_interconnect_0_cam_in_9_s1_readdata                                 : std_logic_vector(31 downto 0); -- cam_in_9:readdata -> mm_interconnect_0:cam_in_9_s1_readdata
	signal mm_interconnect_0_cam_in_9_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:cam_in_9_s1_address -> cam_in_9:address
	signal mm_interconnect_0_cam_in_7_s1_readdata                                 : std_logic_vector(31 downto 0); -- cam_in_7:readdata -> mm_interconnect_0:cam_in_7_s1_readdata
	signal mm_interconnect_0_cam_in_7_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:cam_in_7_s1_address -> cam_in_7:address
	signal mm_interconnect_0_cam_in_6_s1_readdata                                 : std_logic_vector(31 downto 0); -- cam_in_6:readdata -> mm_interconnect_0:cam_in_6_s1_readdata
	signal mm_interconnect_0_cam_in_6_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:cam_in_6_s1_address -> cam_in_6:address
	signal mm_interconnect_0_cam_in_5_s1_readdata                                 : std_logic_vector(31 downto 0); -- cam_in_5:readdata -> mm_interconnect_0:cam_in_5_s1_readdata
	signal mm_interconnect_0_cam_in_5_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:cam_in_5_s1_address -> cam_in_5:address
	signal mm_interconnect_0_cam_in_4_s1_readdata                                 : std_logic_vector(31 downto 0); -- cam_in_4:readdata -> mm_interconnect_0:cam_in_4_s1_readdata
	signal mm_interconnect_0_cam_in_4_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:cam_in_4_s1_address -> cam_in_4:address
	signal mm_interconnect_0_cam_in_3_s1_readdata                                 : std_logic_vector(31 downto 0); -- cam_in_3:readdata -> mm_interconnect_0:cam_in_3_s1_readdata
	signal mm_interconnect_0_cam_in_3_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:cam_in_3_s1_address -> cam_in_3:address
	signal mm_interconnect_0_cam_in_2_s1_readdata                                 : std_logic_vector(31 downto 0); -- cam_in_2:readdata -> mm_interconnect_0:cam_in_2_s1_readdata
	signal mm_interconnect_0_cam_in_2_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:cam_in_2_s1_address -> cam_in_2:address
	signal mm_interconnect_0_cam_in_1_s1_readdata                                 : std_logic_vector(31 downto 0); -- cam_in_1:readdata -> mm_interconnect_0:cam_in_1_s1_readdata
	signal mm_interconnect_0_cam_in_1_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:cam_in_1_s1_address -> cam_in_1:address
	signal mm_interconnect_0_cam_in_0_s1_readdata                                 : std_logic_vector(31 downto 0); -- cam_in_0:readdata -> mm_interconnect_0:cam_in_0_s1_readdata
	signal mm_interconnect_0_cam_in_0_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:cam_in_0_s1_address -> cam_in_0:address
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_chipselect -> JTAG_UART_2nd_Core:av_chipselect
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- JTAG_UART_2nd_Core:av_readdata -> mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest     : std_logic;                     -- JTAG_UART_2nd_Core:av_waitrequest -> mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_address -> JTAG_UART_2nd_Core:av_address
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_writedata -> JTAG_UART_2nd_Core:av_writedata
	signal mm_interconnect_0_nios2_2nd_core_debug_mem_slave_readdata              : std_logic_vector(31 downto 0); -- Nios2_2nd_Core:debug_mem_slave_readdata -> mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_2nd_core_debug_mem_slave_waitrequest           : std_logic;                     -- Nios2_2nd_Core:debug_mem_slave_waitrequest -> mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_2nd_core_debug_mem_slave_debugaccess           : std_logic;                     -- mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_debugaccess -> Nios2_2nd_Core:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_2nd_core_debug_mem_slave_address               : std_logic_vector(8 downto 0);  -- mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_address -> Nios2_2nd_Core:debug_mem_slave_address
	signal mm_interconnect_0_nios2_2nd_core_debug_mem_slave_read                  : std_logic;                     -- mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_read -> Nios2_2nd_Core:debug_mem_slave_read
	signal mm_interconnect_0_nios2_2nd_core_debug_mem_slave_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_byteenable -> Nios2_2nd_Core:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_2nd_core_debug_mem_slave_write                 : std_logic;                     -- mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_write -> Nios2_2nd_Core:debug_mem_slave_write
	signal mm_interconnect_0_nios2_2nd_core_debug_mem_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_writedata -> Nios2_2nd_Core:debug_mem_slave_writedata
	signal irq_mapper_receiver0_irq                                               : std_logic;                     -- JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	signal nios2_irq_irq                                                          : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> Nios2:irq
	signal irq_mapper_001_receiver0_irq                                           : std_logic;                     -- JTAG_UART_2nd_Core:av_irq -> irq_mapper_001:receiver0_irq
	signal nios2_2nd_core_irq_irq                                                 : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> Nios2_2nd_Core:irq
	signal rst_controller_reset_out_reset                                         : std_logic;                     -- rst_controller:reset_out -> [SRAM:reset, mm_interconnect_0:JTAG_UART_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal system_pll_reset_source_reset                                          : std_logic;                     -- System_PLL:reset_source_reset -> [rst_controller:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in2]
	signal rst_controller_001_reset_out_reset                                     : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:Nios2_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal nios2_debug_reset_request_reset                                        : std_logic;                     -- Nios2:debug_reset_request -> [rst_controller_001:reset_in0, rst_controller_003:reset_in1]
	signal rst_controller_002_reset_out_reset                                     : std_logic;                     -- rst_controller_002:reset_out -> [irq_mapper_001:reset, mm_interconnect_0:Nios2_2nd_Core_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal nios2_2nd_core_debug_reset_request_reset                               : std_logic;                     -- Nios2_2nd_Core:debug_reset_request -> [rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal rst_controller_003_reset_out_reset                                     : std_logic;                     -- rst_controller_003:reset_out -> [mm_interconnect_0:cam_in_8_reset_reset_bridge_in_reset_reset, rst_controller_003_reset_out_reset:in]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv           : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> JTAG_UART:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv          : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> JTAG_UART:av_write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                              : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> SDRAM:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> SDRAM:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                             : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> SDRAM:az_wr_n
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read:inv -> JTAG_UART_2nd_Core:av_read_n
	signal mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write:inv -> JTAG_UART_2nd_Core:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                               : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Flash:i_reset_n, JTAG_UART:rst_n, JTAG_UART_2nd_Core:rst_n, SDRAM:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                           : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> Nios2:reset_n
	signal rst_controller_002_reset_out_reset_ports_inv                           : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> Nios2_2nd_Core:reset_n
	signal rst_controller_003_reset_out_reset_ports_inv                           : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> [cam_in_0:reset_n, cam_in_1:reset_n, cam_in_2:reset_n, cam_in_3:reset_n, cam_in_4:reset_n, cam_in_5:reset_n, cam_in_6:reset_n, cam_in_7:reset_n, cam_in_8:reset_n, cam_in_9:reset_n]

begin

	flash : component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface
		generic map (
			FLASH_MEMORY_ADDRESS_WIDTH => 23
		)
		port map (
			i_avalon_chip_select       => mm_interconnect_0_flash_flash_data_chipselect,           --          flash_data.chipselect
			i_avalon_write             => mm_interconnect_0_flash_flash_data_write,                --                    .write
			i_avalon_read              => mm_interconnect_0_flash_flash_data_read,                 --                    .read
			i_avalon_address           => mm_interconnect_0_flash_flash_data_address,              --                    .address
			i_avalon_byteenable        => mm_interconnect_0_flash_flash_data_byteenable,           --                    .byteenable
			i_avalon_writedata         => mm_interconnect_0_flash_flash_data_writedata,            --                    .writedata
			o_avalon_readdata          => mm_interconnect_0_flash_flash_data_readdata,             --                    .readdata
			o_avalon_waitrequest       => mm_interconnect_0_flash_flash_data_waitrequest,          --                    .waitrequest
			i_clock                    => system_pll_sys_clk_clk,                                  --                 clk.clk
			i_reset_n                  => rst_controller_reset_out_reset_ports_inv,                --               reset.reset_n
			FL_ADDR                    => flash_ADDR,                                              --         conduit_end.export
			FL_CE_N                    => flash_CE_N,                                              --                    .export
			FL_OE_N                    => flash_OE_N,                                              --                    .export
			FL_WE_N                    => flash_WE_N,                                              --                    .export
			FL_RST_N                   => flash_RST_N,                                             --                    .export
			FL_DQ                      => flash_DQ,                                                --                    .export
			i_avalon_erase_write       => mm_interconnect_0_flash_flash_erase_control_write,       -- flash_erase_control.write
			i_avalon_erase_read        => mm_interconnect_0_flash_flash_erase_control_read,        --                    .read
			i_avalon_erase_byteenable  => mm_interconnect_0_flash_flash_erase_control_byteenable,  --                    .byteenable
			i_avalon_erase_writedata   => mm_interconnect_0_flash_flash_erase_control_writedata,   --                    .writedata
			i_avalon_erase_chip_select => mm_interconnect_0_flash_flash_erase_control_chipselect,  --                    .chipselect
			o_avalon_erase_readdata    => mm_interconnect_0_flash_flash_erase_control_readdata,    --                    .readdata
			o_avalon_erase_waitrequest => mm_interconnect_0_flash_flash_erase_control_waitrequest  --                    .waitrequest
		);

	jtag_uart : component nios_system_JTAG_UART
		port map (
			clk            => system_pll_sys_clk_clk,                                        --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	jtag_uart_2nd_core : component nios_system_JTAG_UART
		port map (
			clk            => system_pll_sys_clk_clk,                                                 --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                               --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_001_receiver0_irq                                            --               irq.irq
		);

	nios2 : component nios_system_Nios2
		port map (
			clk                                 => system_pll_sys_clk_clk,                              --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,        --                     reset.reset_n
			d_address                           => nios2_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_data_master_read,                              --                          .read
			d_readdata                          => nios2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_data_master_write,                             --                          .write
			d_writedata                         => nios2_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	nios2_2nd_core : component nios_system_Nios2_2nd_Core
		port map (
			clk                                 => system_pll_sys_clk_clk,                                       --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,                 --                     reset.reset_n
			d_address                           => nios2_2nd_core_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_2nd_core_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_2nd_core_data_master_read,                              --                          .read
			d_readdata                          => nios2_2nd_core_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_2nd_core_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_2nd_core_data_master_write,                             --                          .write
			d_writedata                         => nios2_2nd_core_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_2nd_core_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_2nd_core_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_2nd_core_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_2nd_core_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_2nd_core_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_2nd_core_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_2nd_core_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_2nd_core_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                          -- custom_instruction_master.readra
		);

	sdram : component nios_system_SDRAM
		port map (
			clk            => system_pll_sys_clk_clk,                          --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	sram : component nios_system_SRAM
		port map (
			clk           => system_pll_sys_clk_clk,                                 --                clk.clk
			reset         => rst_controller_reset_out_reset,                         --              reset.reset
			SRAM_DQ       => sram_DQ,                                                -- external_interface.export
			SRAM_ADDR     => sram_ADDR,                                              --                   .export
			SRAM_LB_N     => sram_LB_N,                                              --                   .export
			SRAM_UB_N     => sram_UB_N,                                              --                   .export
			SRAM_CE_N     => sram_CE_N,                                              --                   .export
			SRAM_OE_N     => sram_OE_N,                                              --                   .export
			SRAM_WE_N     => sram_WE_N,                                              --                   .export
			address       => mm_interconnect_0_sram_avalon_sram_slave_address,       --  avalon_sram_slave.address
			byteenable    => mm_interconnect_0_sram_avalon_sram_slave_byteenable,    --                   .byteenable
			read          => mm_interconnect_0_sram_avalon_sram_slave_read,          --                   .read
			write         => mm_interconnect_0_sram_avalon_sram_slave_write,         --                   .write
			writedata     => mm_interconnect_0_sram_avalon_sram_slave_writedata,     --                   .writedata
			readdata      => mm_interconnect_0_sram_avalon_sram_slave_readdata,      --                   .readdata
			readdatavalid => mm_interconnect_0_sram_avalon_sram_slave_readdatavalid  --                   .readdatavalid
		);

	system_pll : component nios_system_System_PLL
		port map (
			ref_clk_clk        => system_pll_ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => system_pll_ref_reset_reset,    --    ref_reset.reset
			sys_clk_clk        => system_pll_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                 --    sdram_clk.clk
			reset_source_reset => system_pll_reset_source_reset  -- reset_source.reset
		);

	cam_in_0 : component nios_system_cam_in_0
		port map (
			clk      => system_pll_sys_clk_clk,                       --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_cam_in_0_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_cam_in_0_s1_readdata,       --                    .readdata
			in_port  => cam_in_0_external_connection_export           -- external_connection.export
		);

	cam_in_1 : component nios_system_cam_in_0
		port map (
			clk      => system_pll_sys_clk_clk,                       --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_cam_in_1_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_cam_in_1_s1_readdata,       --                    .readdata
			in_port  => cam_in_1_external_connection_export           -- external_connection.export
		);

	cam_in_2 : component nios_system_cam_in_0
		port map (
			clk      => system_pll_sys_clk_clk,                       --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_cam_in_2_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_cam_in_2_s1_readdata,       --                    .readdata
			in_port  => cam_in_2_external_connection_export           -- external_connection.export
		);

	cam_in_3 : component nios_system_cam_in_0
		port map (
			clk      => system_pll_sys_clk_clk,                       --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_cam_in_3_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_cam_in_3_s1_readdata,       --                    .readdata
			in_port  => cam_in_3_external_connection_export           -- external_connection.export
		);

	cam_in_4 : component nios_system_cam_in_0
		port map (
			clk      => system_pll_sys_clk_clk,                       --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_cam_in_4_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_cam_in_4_s1_readdata,       --                    .readdata
			in_port  => cam_in_4_external_connection_export           -- external_connection.export
		);

	cam_in_5 : component nios_system_cam_in_0
		port map (
			clk      => system_pll_sys_clk_clk,                       --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_cam_in_5_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_cam_in_5_s1_readdata,       --                    .readdata
			in_port  => cam_in_5_external_connection_export           -- external_connection.export
		);

	cam_in_6 : component nios_system_cam_in_0
		port map (
			clk      => system_pll_sys_clk_clk,                       --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_cam_in_6_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_cam_in_6_s1_readdata,       --                    .readdata
			in_port  => cam_in_6_external_connection_export           -- external_connection.export
		);

	cam_in_7 : component nios_system_cam_in_0
		port map (
			clk      => system_pll_sys_clk_clk,                       --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_cam_in_7_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_cam_in_7_s1_readdata,       --                    .readdata
			in_port  => cam_in_7_external_connection_export           -- external_connection.export
		);

	cam_in_8 : component nios_system_cam_in_0
		port map (
			clk      => system_pll_sys_clk_clk,                       --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_cam_in_8_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_cam_in_8_s1_readdata,       --                    .readdata
			in_port  => cam_in_8_external_connection_export           -- external_connection.export
		);

	cam_in_9 : component nios_system_cam_in_0
		port map (
			clk      => system_pll_sys_clk_clk,                       --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_cam_in_9_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_cam_in_9_s1_readdata,       --                    .readdata
			in_port  => cam_in_9_external_connection_export           -- external_connection.export
		);

	mm_interconnect_0 : component nios_system_mm_interconnect_0
		port map (
			System_PLL_sys_clk_clk                           => system_pll_sys_clk_clk,                                             --                         System_PLL_sys_clk.clk
			cam_in_8_reset_reset_bridge_in_reset_reset       => rst_controller_003_reset_out_reset,                                 --       cam_in_8_reset_reset_bridge_in_reset.reset
			JTAG_UART_reset_reset_bridge_in_reset_reset      => rst_controller_reset_out_reset,                                     --      JTAG_UART_reset_reset_bridge_in_reset.reset
			Nios2_2nd_Core_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                                 -- Nios2_2nd_Core_reset_reset_bridge_in_reset.reset
			Nios2_reset_reset_bridge_in_reset_reset          => rst_controller_001_reset_out_reset,                                 --          Nios2_reset_reset_bridge_in_reset.reset
			Nios2_data_master_address                        => nios2_data_master_address,                                          --                          Nios2_data_master.address
			Nios2_data_master_waitrequest                    => nios2_data_master_waitrequest,                                      --                                           .waitrequest
			Nios2_data_master_byteenable                     => nios2_data_master_byteenable,                                       --                                           .byteenable
			Nios2_data_master_read                           => nios2_data_master_read,                                             --                                           .read
			Nios2_data_master_readdata                       => nios2_data_master_readdata,                                         --                                           .readdata
			Nios2_data_master_write                          => nios2_data_master_write,                                            --                                           .write
			Nios2_data_master_writedata                      => nios2_data_master_writedata,                                        --                                           .writedata
			Nios2_data_master_debugaccess                    => nios2_data_master_debugaccess,                                      --                                           .debugaccess
			Nios2_instruction_master_address                 => nios2_instruction_master_address,                                   --                   Nios2_instruction_master.address
			Nios2_instruction_master_waitrequest             => nios2_instruction_master_waitrequest,                               --                                           .waitrequest
			Nios2_instruction_master_read                    => nios2_instruction_master_read,                                      --                                           .read
			Nios2_instruction_master_readdata                => nios2_instruction_master_readdata,                                  --                                           .readdata
			Nios2_instruction_master_readdatavalid           => nios2_instruction_master_readdatavalid,                             --                                           .readdatavalid
			Nios2_2nd_Core_data_master_address               => nios2_2nd_core_data_master_address,                                 --                 Nios2_2nd_Core_data_master.address
			Nios2_2nd_Core_data_master_waitrequest           => nios2_2nd_core_data_master_waitrequest,                             --                                           .waitrequest
			Nios2_2nd_Core_data_master_byteenable            => nios2_2nd_core_data_master_byteenable,                              --                                           .byteenable
			Nios2_2nd_Core_data_master_read                  => nios2_2nd_core_data_master_read,                                    --                                           .read
			Nios2_2nd_Core_data_master_readdata              => nios2_2nd_core_data_master_readdata,                                --                                           .readdata
			Nios2_2nd_Core_data_master_write                 => nios2_2nd_core_data_master_write,                                   --                                           .write
			Nios2_2nd_Core_data_master_writedata             => nios2_2nd_core_data_master_writedata,                               --                                           .writedata
			Nios2_2nd_Core_data_master_debugaccess           => nios2_2nd_core_data_master_debugaccess,                             --                                           .debugaccess
			Nios2_2nd_Core_instruction_master_address        => nios2_2nd_core_instruction_master_address,                          --          Nios2_2nd_Core_instruction_master.address
			Nios2_2nd_Core_instruction_master_waitrequest    => nios2_2nd_core_instruction_master_waitrequest,                      --                                           .waitrequest
			Nios2_2nd_Core_instruction_master_read           => nios2_2nd_core_instruction_master_read,                             --                                           .read
			Nios2_2nd_Core_instruction_master_readdata       => nios2_2nd_core_instruction_master_readdata,                         --                                           .readdata
			Nios2_2nd_Core_instruction_master_readdatavalid  => nios2_2nd_core_instruction_master_readdatavalid,                    --                                           .readdatavalid
			cam_in_0_s1_address                              => mm_interconnect_0_cam_in_0_s1_address,                              --                                cam_in_0_s1.address
			cam_in_0_s1_readdata                             => mm_interconnect_0_cam_in_0_s1_readdata,                             --                                           .readdata
			cam_in_1_s1_address                              => mm_interconnect_0_cam_in_1_s1_address,                              --                                cam_in_1_s1.address
			cam_in_1_s1_readdata                             => mm_interconnect_0_cam_in_1_s1_readdata,                             --                                           .readdata
			cam_in_2_s1_address                              => mm_interconnect_0_cam_in_2_s1_address,                              --                                cam_in_2_s1.address
			cam_in_2_s1_readdata                             => mm_interconnect_0_cam_in_2_s1_readdata,                             --                                           .readdata
			cam_in_3_s1_address                              => mm_interconnect_0_cam_in_3_s1_address,                              --                                cam_in_3_s1.address
			cam_in_3_s1_readdata                             => mm_interconnect_0_cam_in_3_s1_readdata,                             --                                           .readdata
			cam_in_4_s1_address                              => mm_interconnect_0_cam_in_4_s1_address,                              --                                cam_in_4_s1.address
			cam_in_4_s1_readdata                             => mm_interconnect_0_cam_in_4_s1_readdata,                             --                                           .readdata
			cam_in_5_s1_address                              => mm_interconnect_0_cam_in_5_s1_address,                              --                                cam_in_5_s1.address
			cam_in_5_s1_readdata                             => mm_interconnect_0_cam_in_5_s1_readdata,                             --                                           .readdata
			cam_in_6_s1_address                              => mm_interconnect_0_cam_in_6_s1_address,                              --                                cam_in_6_s1.address
			cam_in_6_s1_readdata                             => mm_interconnect_0_cam_in_6_s1_readdata,                             --                                           .readdata
			cam_in_7_s1_address                              => mm_interconnect_0_cam_in_7_s1_address,                              --                                cam_in_7_s1.address
			cam_in_7_s1_readdata                             => mm_interconnect_0_cam_in_7_s1_readdata,                             --                                           .readdata
			cam_in_8_s1_address                              => mm_interconnect_0_cam_in_8_s1_address,                              --                                cam_in_8_s1.address
			cam_in_8_s1_readdata                             => mm_interconnect_0_cam_in_8_s1_readdata,                             --                                           .readdata
			cam_in_9_s1_address                              => mm_interconnect_0_cam_in_9_s1_address,                              --                                cam_in_9_s1.address
			cam_in_9_s1_readdata                             => mm_interconnect_0_cam_in_9_s1_readdata,                             --                                           .readdata
			Flash_flash_data_address                         => mm_interconnect_0_flash_flash_data_address,                         --                           Flash_flash_data.address
			Flash_flash_data_write                           => mm_interconnect_0_flash_flash_data_write,                           --                                           .write
			Flash_flash_data_read                            => mm_interconnect_0_flash_flash_data_read,                            --                                           .read
			Flash_flash_data_readdata                        => mm_interconnect_0_flash_flash_data_readdata,                        --                                           .readdata
			Flash_flash_data_writedata                       => mm_interconnect_0_flash_flash_data_writedata,                       --                                           .writedata
			Flash_flash_data_byteenable                      => mm_interconnect_0_flash_flash_data_byteenable,                      --                                           .byteenable
			Flash_flash_data_waitrequest                     => mm_interconnect_0_flash_flash_data_waitrequest,                     --                                           .waitrequest
			Flash_flash_data_chipselect                      => mm_interconnect_0_flash_flash_data_chipselect,                      --                                           .chipselect
			Flash_flash_erase_control_write                  => mm_interconnect_0_flash_flash_erase_control_write,                  --                  Flash_flash_erase_control.write
			Flash_flash_erase_control_read                   => mm_interconnect_0_flash_flash_erase_control_read,                   --                                           .read
			Flash_flash_erase_control_readdata               => mm_interconnect_0_flash_flash_erase_control_readdata,               --                                           .readdata
			Flash_flash_erase_control_writedata              => mm_interconnect_0_flash_flash_erase_control_writedata,              --                                           .writedata
			Flash_flash_erase_control_byteenable             => mm_interconnect_0_flash_flash_erase_control_byteenable,             --                                           .byteenable
			Flash_flash_erase_control_waitrequest            => mm_interconnect_0_flash_flash_erase_control_waitrequest,            --                                           .waitrequest
			Flash_flash_erase_control_chipselect             => mm_interconnect_0_flash_flash_erase_control_chipselect,             --                                           .chipselect
			JTAG_UART_avalon_jtag_slave_address              => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,              --                JTAG_UART_avalon_jtag_slave.address
			JTAG_UART_avalon_jtag_slave_write                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,                --                                           .write
			JTAG_UART_avalon_jtag_slave_read                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                 --                                           .read
			JTAG_UART_avalon_jtag_slave_readdata             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,             --                                           .readdata
			JTAG_UART_avalon_jtag_slave_writedata            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,            --                                           .writedata
			JTAG_UART_avalon_jtag_slave_waitrequest          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,          --                                           .waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,           --                                           .chipselect
			JTAG_UART_2nd_Core_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address,     --       JTAG_UART_2nd_Core_avalon_jtag_slave.address
			JTAG_UART_2nd_Core_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write,       --                                           .write
			JTAG_UART_2nd_Core_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read,        --                                           .read
			JTAG_UART_2nd_Core_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata,    --                                           .readdata
			JTAG_UART_2nd_Core_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata,   --                                           .writedata
			JTAG_UART_2nd_Core_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest, --                                           .waitrequest
			JTAG_UART_2nd_Core_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect,  --                                           .chipselect
			Nios2_debug_mem_slave_address                    => mm_interconnect_0_nios2_debug_mem_slave_address,                    --                      Nios2_debug_mem_slave.address
			Nios2_debug_mem_slave_write                      => mm_interconnect_0_nios2_debug_mem_slave_write,                      --                                           .write
			Nios2_debug_mem_slave_read                       => mm_interconnect_0_nios2_debug_mem_slave_read,                       --                                           .read
			Nios2_debug_mem_slave_readdata                   => mm_interconnect_0_nios2_debug_mem_slave_readdata,                   --                                           .readdata
			Nios2_debug_mem_slave_writedata                  => mm_interconnect_0_nios2_debug_mem_slave_writedata,                  --                                           .writedata
			Nios2_debug_mem_slave_byteenable                 => mm_interconnect_0_nios2_debug_mem_slave_byteenable,                 --                                           .byteenable
			Nios2_debug_mem_slave_waitrequest                => mm_interconnect_0_nios2_debug_mem_slave_waitrequest,                --                                           .waitrequest
			Nios2_debug_mem_slave_debugaccess                => mm_interconnect_0_nios2_debug_mem_slave_debugaccess,                --                                           .debugaccess
			Nios2_2nd_Core_debug_mem_slave_address           => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_address,           --             Nios2_2nd_Core_debug_mem_slave.address
			Nios2_2nd_Core_debug_mem_slave_write             => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_write,             --                                           .write
			Nios2_2nd_Core_debug_mem_slave_read              => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_read,              --                                           .read
			Nios2_2nd_Core_debug_mem_slave_readdata          => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_readdata,          --                                           .readdata
			Nios2_2nd_Core_debug_mem_slave_writedata         => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_writedata,         --                                           .writedata
			Nios2_2nd_Core_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_byteenable,        --                                           .byteenable
			Nios2_2nd_Core_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_waitrequest,       --                                           .waitrequest
			Nios2_2nd_Core_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_2nd_core_debug_mem_slave_debugaccess,       --                                           .debugaccess
			SDRAM_s1_address                                 => mm_interconnect_0_sdram_s1_address,                                 --                                   SDRAM_s1.address
			SDRAM_s1_write                                   => mm_interconnect_0_sdram_s1_write,                                   --                                           .write
			SDRAM_s1_read                                    => mm_interconnect_0_sdram_s1_read,                                    --                                           .read
			SDRAM_s1_readdata                                => mm_interconnect_0_sdram_s1_readdata,                                --                                           .readdata
			SDRAM_s1_writedata                               => mm_interconnect_0_sdram_s1_writedata,                               --                                           .writedata
			SDRAM_s1_byteenable                              => mm_interconnect_0_sdram_s1_byteenable,                              --                                           .byteenable
			SDRAM_s1_readdatavalid                           => mm_interconnect_0_sdram_s1_readdatavalid,                           --                                           .readdatavalid
			SDRAM_s1_waitrequest                             => mm_interconnect_0_sdram_s1_waitrequest,                             --                                           .waitrequest
			SDRAM_s1_chipselect                              => mm_interconnect_0_sdram_s1_chipselect,                              --                                           .chipselect
			SRAM_avalon_sram_slave_address                   => mm_interconnect_0_sram_avalon_sram_slave_address,                   --                     SRAM_avalon_sram_slave.address
			SRAM_avalon_sram_slave_write                     => mm_interconnect_0_sram_avalon_sram_slave_write,                     --                                           .write
			SRAM_avalon_sram_slave_read                      => mm_interconnect_0_sram_avalon_sram_slave_read,                      --                                           .read
			SRAM_avalon_sram_slave_readdata                  => mm_interconnect_0_sram_avalon_sram_slave_readdata,                  --                                           .readdata
			SRAM_avalon_sram_slave_writedata                 => mm_interconnect_0_sram_avalon_sram_slave_writedata,                 --                                           .writedata
			SRAM_avalon_sram_slave_byteenable                => mm_interconnect_0_sram_avalon_sram_slave_byteenable,                --                                           .byteenable
			SRAM_avalon_sram_slave_readdatavalid             => mm_interconnect_0_sram_avalon_sram_slave_readdatavalid              --                                           .readdatavalid
		);

	irq_mapper : component nios_system_irq_mapper
		port map (
			clk           => system_pll_sys_clk_clk,             --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			sender_irq    => nios2_irq_irq                       --    sender.irq
		);

	irq_mapper_001 : component nios_system_irq_mapper
		port map (
			clk           => system_pll_sys_clk_clk,             --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios2_2nd_core_irq_irq              --    sender.irq
		);

	rst_controller : component nios_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => system_pll_reset_source_reset,  -- reset_in0.reset
			clk            => system_pll_sys_clk_clk,         --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component nios_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_debug_reset_request_reset,    -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,      -- reset_in1.reset
			clk            => system_pll_sys_clk_clk,             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component nios_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_2nd_core_debug_reset_request_reset, -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,            -- reset_in1.reset
			clk            => system_pll_sys_clk_clk,                   --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,       -- reset_out.reset
			reset_req      => open,                                     -- (terminated)
			reset_req_in0  => '0',                                      -- (terminated)
			reset_req_in1  => '0',                                      -- (terminated)
			reset_in2      => '0',                                      -- (terminated)
			reset_req_in2  => '0',                                      -- (terminated)
			reset_in3      => '0',                                      -- (terminated)
			reset_req_in3  => '0',                                      -- (terminated)
			reset_in4      => '0',                                      -- (terminated)
			reset_req_in4  => '0',                                      -- (terminated)
			reset_in5      => '0',                                      -- (terminated)
			reset_req_in5  => '0',                                      -- (terminated)
			reset_in6      => '0',                                      -- (terminated)
			reset_req_in6  => '0',                                      -- (terminated)
			reset_in7      => '0',                                      -- (terminated)
			reset_req_in7  => '0',                                      -- (terminated)
			reset_in8      => '0',                                      -- (terminated)
			reset_req_in8  => '0',                                      -- (terminated)
			reset_in9      => '0',                                      -- (terminated)
			reset_req_in9  => '0',                                      -- (terminated)
			reset_in10     => '0',                                      -- (terminated)
			reset_req_in10 => '0',                                      -- (terminated)
			reset_in11     => '0',                                      -- (terminated)
			reset_req_in11 => '0',                                      -- (terminated)
			reset_in12     => '0',                                      -- (terminated)
			reset_req_in12 => '0',                                      -- (terminated)
			reset_in13     => '0',                                      -- (terminated)
			reset_req_in13 => '0',                                      -- (terminated)
			reset_in14     => '0',                                      -- (terminated)
			reset_req_in14 => '0',                                      -- (terminated)
			reset_in15     => '0',                                      -- (terminated)
			reset_req_in15 => '0'                                       -- (terminated)
		);

	rst_controller_003 : component nios_system_rst_controller_003
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_2nd_core_debug_reset_request_reset, -- reset_in0.reset
			reset_in1      => nios2_debug_reset_request_reset,          -- reset_in1.reset
			reset_in2      => system_pll_reset_source_reset,            -- reset_in2.reset
			clk            => system_pll_sys_clk_clk,                   --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,       -- reset_out.reset
			reset_req      => open,                                     -- (terminated)
			reset_req_in0  => '0',                                      -- (terminated)
			reset_req_in1  => '0',                                      -- (terminated)
			reset_req_in2  => '0',                                      -- (terminated)
			reset_in3      => '0',                                      -- (terminated)
			reset_req_in3  => '0',                                      -- (terminated)
			reset_in4      => '0',                                      -- (terminated)
			reset_req_in4  => '0',                                      -- (terminated)
			reset_in5      => '0',                                      -- (terminated)
			reset_req_in5  => '0',                                      -- (terminated)
			reset_in6      => '0',                                      -- (terminated)
			reset_req_in6  => '0',                                      -- (terminated)
			reset_in7      => '0',                                      -- (terminated)
			reset_req_in7  => '0',                                      -- (terminated)
			reset_in8      => '0',                                      -- (terminated)
			reset_req_in8  => '0',                                      -- (terminated)
			reset_in9      => '0',                                      -- (terminated)
			reset_req_in9  => '0',                                      -- (terminated)
			reset_in10     => '0',                                      -- (terminated)
			reset_req_in10 => '0',                                      -- (terminated)
			reset_in11     => '0',                                      -- (terminated)
			reset_req_in11 => '0',                                      -- (terminated)
			reset_in12     => '0',                                      -- (terminated)
			reset_req_in12 => '0',                                      -- (terminated)
			reset_in13     => '0',                                      -- (terminated)
			reset_req_in13 => '0',                                      -- (terminated)
			reset_in14     => '0',                                      -- (terminated)
			reset_req_in14 => '0',                                      -- (terminated)
			reset_in15     => '0',                                      -- (terminated)
			reset_req_in15 => '0'                                       -- (terminated)
		);

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

end architecture rtl; -- of nios_system
