--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.numeric_std.all;
--
--entity Colour_Recognition_register is
--  Port (
--    activated			: in std_logic;
--    clk_i 				: in std_logic;
--	 dpixel 				: in std_logic_vector (11 downto 0);
--    address_second 	: in std_logic_vector (16 downto 0);
--	 colour				: out std_logic_vector (11 downto 0);
--	 pixel				: out std_logic_vector (11 downto 0);
--	 
--	 -- here we placed all the variables that will be used by the C code
--	 -- empty: 				001
--	 -- friendly stone:	010
--	 -- friendly king:	011
--	 -- enemy stone:		100
--	 -- enemy king:		101
--	 vak_1 				: out std_logic_vector(2 downto 0);
--	 vak_2 				: out std_logic_vector(2 downto 0);
--	 vak_3 				: out std_logic_vector(2 downto 0);
--	 vak_4 				: out std_logic_vector(2 downto 0);
--	 vak_5 				: out std_logic_vector(2 downto 0);
--	 vak_6 				: out std_logic_vector(2 downto 0);
--	 vak_7 				: out std_logic_vector(2 downto 0);
--	 vak_8 				: out std_logic_vector(2 downto 0);
--	 vak_9 				: out std_logic_vector(2 downto 0);
--	 vak_10 				: out std_logic_vector(2 downto 0);
--	 vak_11 				: out std_logic_vector(2 downto 0);
--	 vak_12 				: out std_logic_vector(2 downto 0);
--	 vak_13 				: out std_logic_vector(2 downto 0);
--	 vak_14 				: out std_logic_vector(2 downto 0);
--	 vak_15				: out std_logic_vector(2 downto 0);
--	 vak_16 				: out std_logic_vector(2 downto 0);
--	 vak_17 				: out std_logic_vector(2 downto 0);
--	 vak_18 				: out std_logic_vector(2 downto 0);
--	 vak_19 				: out std_logic_vector(2 downto 0);
--	 vak_20 				: out std_logic_vector(2 downto 0);
--	 vak_21 				: out std_logic_vector(2 downto 0);
--	 vak_22 				: out std_logic_vector(2 downto 0);
--	 vak_23 				: out std_logic_vector(2 downto 0);
--	 vak_24 				: out std_logic_vector(2 downto 0);
--	 vak_25 				: out std_logic_vector(2 downto 0);
--	 vak_26 				: out std_logic_vector(2 downto 0);
--	 vak_27 				: out std_logic_vector(2 downto 0);
--	 vak_28 				: out std_logic_vector(2 downto 0);
--	 vak_29 				: out std_logic_vector(2 downto 0);
--	 vak_30 				: out std_logic_vector(2 downto 0);
--	 vak_31 				: out std_logic_vector(2 downto 0);
--	 vak_32 				: out std_logic_vector(2 downto 0);
--	 vak_33 				: out std_logic_vector(2 downto 0);
--	 vak_34 				: out std_logic_vector(2 downto 0);
--	 vak_35 				: out std_logic_vector(2 downto 0);
--	 vak_36 				: out std_logic_vector(2 downto 0);
--	 vak_37 				: out std_logic_vector(2 downto 0);
--	 vak_38 				: out std_logic_vector(2 downto 0);
--	 vak_39 				: out std_logic_vector(2 downto 0);
--	 vak_40 				: out std_logic_vector(2 downto 0);
--	 vak_41 				: out std_logic_vector(2 downto 0);
--	 vak_42 				: out std_logic_vector(2 downto 0);
--	 vak_43 				: out std_logic_vector(2 downto 0);
--	 vak_44 				: out std_logic_vector(2 downto 0);
--	 vak_45 				: out std_logic_vector(2 downto 0);
--	 vak_46 				: out std_logic_vector(2 downto 0);
--	 vak_47 				: out std_logic_vector(2 downto 0);
--	 vak_48 				: out std_logic_vector(2 downto 0);
--	 vak_49 				: out std_logic_vector(2 downto 0);
--	 vak_50 				: out std_logic_vector(2 downto 0)
--  );  
--end Colour_Recognition_register;
--
--architecture Recognize of Colour_Recognition is
--
----signal red					: unsigned(7 downto 0);				-- bevat het totaal aantal rood van een vakje
----signal green				: unsigned(7 downto 0);				-- bevat het totaal aantal groen van een vakje
----signal blue					: unsigned(7 downto 0);				-- bevat het totaal aantal blauw van een vakje
----signal temp_red			: unsigned(3 downto 0);				-- bevat van 1 pixel de kleur rood
----signal temp_green			: unsigned(3 downto 0);				-- bevat van 1 pixel de kleur groen
----signal temp_blue			: unsigned(3 downto 0);				-- bevat van 1 pixel de kleur blauw
----signal temp_address		: unsigned(16 downto 0);			-- bevat de unsigned versie van het address
--signal frameCounter		: std_logic_vector(1 downto 0);	-- bevat hoe vaak er een frame is gebruikt per knop indruk. 00: 0 frames, 01: 1 frame, 10: meer dan 1 frame
--  
--  type redArray is array (0 to 49) of unsigned(5 downto 0);
--  signal red : redArray;
--  type greenArray is array (0 to 49) of unsigned(5 downto 0);
--  signal green : greenArray;
--  type blueArray is array (0 to 49) of unsigned(5 downto 0);
--  signal blue : blueArray;
--  
----  type temp_redArray is array (0 to 49) of unsigned(3 downto 0);
----  signal temp_red : temp_redArray;
----  type temp_greenArray is array (0 to 49) of unsigned(3 downto 0);
----  signal temp_green : temp_greenArray;
----  type temp_blueArray is array (0 to 49) of unsigned(3 downto 0);
----  signal temp_blue : temp_blueArray;
--  
--  -- array die de addressen van de vakjes bevat waar er kleur herkenning moet uitgevoerd worden
--  -- (vak nummer)(addres van de pixel links boven van het vak)
--  type limitPixelArray is array (0 to 49) of unsigned(16 downto 0);
--  signal limitPixel_main : limitPixelArray;
--  
--  -- array die bevat wat een vakje nou eigenlijk bevat. friendly, enemy, ....
--  -- (vak nummer)(inhoud)
--  type vakInhoudArray is array (0 to 49) of std_logic_vector(2 downto 0);
--  signal vakInhoud_main : vakInhoudArray;
--  
--  -- array die de pixel bevat die uiteindelijk terug naar de vga gaat
--  -- in essentie zouden al deze waardes hetzelfde moeten zijn
--  -- (vaknummer)(pixel)
--  type pixelArray is array (0 to 49) of std_logic_vector(11 downto 0);
--  signal pixel_main : pixelArray;
--  
--  -- array die de gemiddelde kleur bevat van een vakje
--  -- (vaknummer)(kleur)
--  type colourArray is array (0 to 49) of std_logic_vector(11 downto 0);
--  signal colour_main : colourArray;
--  
--  signal activeSend 		: std_logic := '0';
--  signal activeInhoud 	: std_logic := '0';
--  
--  signal limitPixel		: unsigned(16 downto 0);
--  
--  signal number			: integer range 0 to 49;
--
--begin
--	limitPixel <= to_unsigned(752, 17);
--	
--	-- hier worden alle addressen opgeslagen van de pixel die links boven in een vakje zit
--	-- eerst werd dit met een functie gedaan, alleen bleek dit zeer inefficient te zijn
--	limitPixel_main(0) <= to_unsigned(752, 17);
--	limitPixel_main(1) <= to_unsigned(784, 17);
--	limitPixel_main(2) <= to_unsigned(816, 17);
--	limitPixel_main(3) <= to_unsigned(848, 17);
--	limitPixel_main(4) <= to_unsigned(880, 17);
--	limitPixel_main(5) <= to_unsigned(5856, 17);
--	limitPixel_main(6) <= to_unsigned(5888, 17);
--	limitPixel_main(7) <= to_unsigned(5920, 17);
--	limitPixel_main(8) <= to_unsigned(5952, 17);
--	limitPixel_main(9) <= to_unsigned(5984, 17);
--	limitPixel_main(10) <= to_unsigned(10992, 17);
--	limitPixel_main(11) <= to_unsigned(11024, 17);
--	limitPixel_main(12) <= to_unsigned(11056, 17);
--	limitPixel_main(13) <= to_unsigned(11088, 17);
--	limitPixel_main(14) <= to_unsigned(11120, 17);
--	limitPixel_main(15) <= to_unsigned(16096, 17);
--	limitPixel_main(16) <= to_unsigned(16128, 17);
--	limitPixel_main(17) <= to_unsigned(16160, 17);
--	limitPixel_main(18) <= to_unsigned(16192, 17);
--	limitPixel_main(19) <= to_unsigned(16224, 17);
--	limitPixel_main(20) <= to_unsigned(21232, 17);
--	limitPixel_main(21) <= to_unsigned(21264, 17);
--	limitPixel_main(22) <= to_unsigned(21296, 17);
--	limitPixel_main(23) <= to_unsigned(21328, 17);
--	limitPixel_main(24) <= to_unsigned(21360, 17);
--	limitPixel_main(25) <= to_unsigned(26336, 17);
--	limitPixel_main(26) <= to_unsigned(26368, 17);
--	limitPixel_main(27) <= to_unsigned(26400, 17);
--	limitPixel_main(28) <= to_unsigned(26432, 17);
--	limitPixel_main(29) <= to_unsigned(26464, 17);
--	limitPixel_main(30) <= to_unsigned(31472, 17);
--	limitPixel_main(31) <= to_unsigned(31504, 17);
--	limitPixel_main(32) <= to_unsigned(31536, 17);
--	limitPixel_main(33) <= to_unsigned(31568, 17);
--	limitPixel_main(34) <= to_unsigned(31600, 17);
--	limitPixel_main(35) <= to_unsigned(36576, 17);
--	limitPixel_main(36) <= to_unsigned(36608, 17);
--	limitPixel_main(37) <= to_unsigned(36640, 17);
--	limitPixel_main(38) <= to_unsigned(36672, 17);
--	limitPixel_main(39) <= to_unsigned(36704, 17);
--	limitPixel_main(40) <= to_unsigned(41712, 17);
--	limitPixel_main(41) <= to_unsigned(41744, 17);
--	limitPixel_main(42) <= to_unsigned(41776, 17);
--	limitPixel_main(43) <= to_unsigned(41808, 17);
--	limitPixel_main(44) <= to_unsigned(41840, 17);
--	limitPixel_main(45) <= to_unsigned(46816, 17);
--	limitPixel_main(46) <= to_unsigned(46848, 17);
--	limitPixel_main(47) <= to_unsigned(46880, 17);
--	limitPixel_main(48) <= to_unsigned(46912, 17);
--	limitPixel_main(49) <= to_unsigned(46944, 17);
--	
--	process (clk_ii)
--	begin
--		if rising_edge (clk_ii) then
--			pixel <= dapixel;
--			temp_address <= unsigned(address);
--			
--			if (temp_address > (limitPixel_main(49)+960)) then
--				if (temp_address < )limitPixel_main(49)+965)) then
--					number <= 49;
--					go <= '1';
--				end if;
--			end if;
--			if (temp_address > (limitPixel_main(49)+640)) then
--				if (temp_address < )limitPixel_main(49)+645)) then
--					number <= 49;
--					go <= '1';
--				end if;
--			end if;
--			if (temp_address > (limitPixel_main(49)+320)) then
--				if (temp_address < )limitPixel_main(49)+325)) then
--					number <= 49;
--					go <= '1';
--				end if;
--			end if;
--			if (temp_address > (limitPixel_main(49))) then
--				if (temp_address < )limitPixel_main(49)+5)) then
--					number <= 49;
--					go <= '1';
--				end if;
--			end if;
--			
--			if (go = '1') then
--				temp_red <= unsigned(dapixel(11 downto 8));
--				temp_green <= unsigned(dapixel(7 downto 4));
--				temp_blue <= unsigned(dapixel(3 downto 0));
--				red(number) <= red(number) + temp_red;
--				green(number) <= green(number) + temp_green;
--				blue(number) <= blue(number) + temp_green;
--				pixel <= "000011110000";
--				go <= '0';
--			else
--				pixel <= dapixel;
--			end if;
--				if (temp_address = 76799) then
--					if (frameCounter = "01") then
--						for I in 0 to 49 loop
--							colour(I)(11 downto 8) <= std_logic_vector(red(I)(5 downto 2));
--							colour(I)(7 downto 4) <= std_logic_vector(green(I)(5 downto 2));
--							colour(I)(3 downto 0) <= std_logic_vector(blue(I)(5 downto 2));
----							colour <= std_logic_vector(unsigned(dapixel));
--							red <= "00000000";
--							green <= "00000000";
--							blue <= "00000000";
--							frameCounter <= "10";
--						end loop;
--					elsif (frameCounter ="00") then
--						frameCounter <= "01";
--					end if;
--				end if;
--				temp_red <= "0000";
--				temp_green <= "0000";
--				temp_blue <= "0000";
--			else
--				frameCounter <= "00";
--				pixel <= dapixel;
--			end if;
--		end if;
--	end process;
--end Recognize;